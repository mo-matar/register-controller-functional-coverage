// This file is no longer used - scoreboard moved to scoreboard.sv
// TestRegistry moved to test_registry.sv