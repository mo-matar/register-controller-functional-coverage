// Top-level testbench file that includes all components
`include "interface.sv"
`include "reg_ctrl_pkg.sv"
`include "../tests/basic_test.sv"
`include "reg_ctrl_tb.sv"
